module uc_interface(
	
    );


endmodule
